module stopwatch_base(
    input clk, rst,
    output [5:0] seconds_ones_counter;
    output [3:0] seconds_tens_counter;
    output [3:0] minutes_ones_counter;
    output [3:0] minutes_tens_counter;
);
    
endmodule
